library verilog;
use verilog.vl_types.all;
entity dut_if is
end dut_if;
