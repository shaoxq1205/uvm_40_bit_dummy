// `timescale 1 ns / 1 ns
// //Test added by Xiaoqiang
// interface dut_if();
// 	logic clk, rst;
// 	logic [39:0] data_in;
// 	logic [39:0] data_out;

// endinterface